class ethmac_ref;

task run();
	$display("ethmac_ref::run");
endtask

endclass
