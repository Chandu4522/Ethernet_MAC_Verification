class ethmac_ckr;

task run();
	$display("ethmac_ckr::run");
endtask

endclass
