class mii_agent extends uvm_agent;
`uvm_component_utils(mii_agent)
`NEW_COMP

function void build_phase(uvm_phase phase);
	super.build_phase(phase);
endfunction

endclass